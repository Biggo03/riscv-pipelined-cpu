//////////////////////////////////////////////
//                reg_write                 //
//////////////////////////////////////////////
`define WRITE_REG       1'b1
`define NO_WRITE_REG    1'b0

//////////////////////////////////////////////
//                  imm_src                 //
//////////////////////////////////////////////
`define I_EXT           3'b000
`define S_EXT           3'b001
`define B_EXT           3'b010
`define J_EXT           3'b011
`define U_EXT           3'b100
`define CSR_EXT         3'b101
`define NA_EXT          3'b000  // fallback

//////////////////////////////////////////////
//                 alu_src                  //
//////////////////////////////////////////////
`define ALU_SRC_WD      1'b0
`define ALU_SRC_IMM     1'b1
`define ALU_SRC_NA      1'b0    // fallback

//////////////////////////////////////////////
//                mem_write                 //
//////////////////////////////////////////////
`define WRITE_MEM       1'b1
`define NO_WRITE_MEM    1'b0

//////////////////////////////////////////////
//               result_src                 //
//////////////////////////////////////////////
`define RESULT_ALU      3'b000
`define RESULT_PCTARGET 3'b001
`define RESULT_PCPLUS4  3'b010
`define RESULT_IMM_EXT  3'b011
`define RESULT_MEM_DATA 3'b100
`define RESULT_CSR      3'b101
`define RESULT_NA       3'b000   // fallback

//////////////////////////////////////////////
//                branch_op                 //
//////////////////////////////////////////////
`define NON_BRANCH      2'b00
`define JUMP            2'b01
`define BRANCH          2'b11

//////////////////////////////////////////////
//                 width_op                 //
//////////////////////////////////////////////
`define WIDTH_CONST     1'b0
`define WIDTH_PROCESS   1'b1

//////////////////////////////////////////////
//                  alu_op                  //
//////////////////////////////////////////////
`define ALU_OP_ADD      2'b00
`define ALU_OP_SUB      2'b01
`define ALU_OP_PROCESS  2'b10
`define ALU_OP_NA       2'b00 // fallback

//////////////////////////////////////////////
//               alu_control                //
//////////////////////////////////////////////
`define ALU_SRL         4'b0000
`define ALU_SRA         4'b0001
`define ALU_AND         4'b0010
`define ALU_OR          4'b0011
`define ALU_XOR         4'b0100
`define ALU_SLT         4'b0101
`define ALU_SLTU        4'b0110
`define ALU_SLL         4'b0111
`define ALU_ADD         4'b1000
`define ALU_SUB         4'b1001

//////////////////////////////////////////////
//                width_src                 //
//////////////////////////////////////////////
`define WIDTH_32        3'b000
`define WIDTH_16S       3'b010
`define WIDTH_16U       3'b110
`define WIDTH_8S        3'b001
`define WIDTH_8U        3'b101

//////////////////////////////////////////////
//                pc_src                    //
//////////////////////////////////////////////
`define PC_SRC_SEQ_F        2'b00
`define PC_SRC_PRED_F       2'b01
`define PC_SRC_SEQ_E        2'b10
`define PC_SRC_TARGET_E     2'b11

//////////////////////////////////////////////
//             pc_base_src                  //
//////////////////////////////////////////////
`define PC_BASE_PC      1'b0
`define PC_BASE_SRCA    1'b1
`define PC_BASE_NA      1'b0 // fallback

//////////////////////////////////////////////
//                  forward                 //
//////////////////////////////////////////////
`define NO_FORWARD      2'b00
`define WB_FORWARD      2'b01
`define MEM_FORWARD     2'b10

//////////////////////////////////////////////
//                 csr_we                   //
//////////////////////////////////////////////
`define WRITE_CSR       1'b1
`define NO_WRITE_CSR    1'b0

//////////////////////////////////////////////
//               csr_control                //
//////////////////////////////////////////////
`define CSR_PASS        2'b01
`define CSR_SET         2'b10
`define CSR_CLEAR       2'b11
`define CSR_NA          2'b01 // fallback

//////////////////////////////////////////////
//                  csr_src                 //
//////////////////////////////////////////////
`define CSR_SRC_REG         1'b0
`define CSR_SRC_IMM         1'b1
`define CSR_SRC_NA          1'b1 // fallback
