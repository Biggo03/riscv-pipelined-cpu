`timescale 1ns / 1ps
//==============================================================//
//  Module:       memory_stage
//  File:         memory_stage.sv
//  Description:  All logic contained within the memory pipeline stage and it's pipeline register
//
//  Author:       Viggo Wozniak
//  Project:      RISC-V Processor
//  Repository:   https://github.com/Biggo03/RISC-V-Pipelined
//
//  Parameters:   N/A
//
//  Notes:        N/A
//==============================================================//
`include "control_macros.sv"

module memory_stage (
    // Clock & reset_i
    input  logic        clk_i,
    input  logic        reset_i,

    // data inputs
    input  logic [31:0] instr_e_i,
    input  logic [31:0] alu_result_e_i,
    input  logic [31:0] write_data_e_i,
    input  logic [31:0] pc_target_e_i,
    input  logic [31:0] pc_plus4_e_i,
    input  logic [31:0] imm_ext_e_i,
    input  logic [31:0] read_data_m_i,
    input  logic [31:0] csr_result_e_i,
    input  logic [31:0] csr_data_e_i,
    input  logic [11:0] csr_addr_e_i,
    input  logic [4:0]  rd_e_i,

    // Control inputs
    input  logic        valid_e_i,
    input  logic [2:0]  width_src_e_i,
    input  logic [2:0]  result_src_e_i,
    input  logic        mem_write_e_i,
    input  logic        reg_write_e_i,
    input  logic        csr_we_e_i,
    input  logic        stall_m_i,

    // data outputs
    output logic [31:0] instr_m_o,
    output logic [31:0] reduced_data_m_o,
    output logic [31:0] alu_result_m_o,
    output logic [31:0] write_data_m_o,
    output logic [31:0] pc_target_m_o,
    output logic [31:0] pc_plus4_m_o,
    output logic [31:0] imm_ext_m_o,
    output logic [31:0] forward_data_m_o,
    output logic [31:0] csr_result_m_o,
    output logic [31:0] csr_data_m_o,
    output logic [11:0] csr_addr_m_o,
    output logic [4:0]  rd_m_o,

    // Control outputs
    output logic        valid_m_o,
    output logic [2:0]  result_src_m_o,
    output logic [2:0]  width_src_m_o,
    output logic        mem_write_m_o,
    output logic        reg_write_m_o,
    output logic        csr_we_m_o
);

    // ----- Pipeline data type -----
    typedef struct packed {
        logic [31:0] instr;
        logic        valid;
        logic [31:0] alu_result;
        logic [31:0] write_data;
        logic [31:0] pc_target;
        logic [31:0] pc_plus4;
        logic [31:0] imm_ext;
        logic [31:0] csr_result;
        logic [31:0] csr_data;
        logic [11:0] csr_addr;
        logic [4:0]  rd;
        logic [2:0]  width_src;
        logic [2:0]  result_src;
        logic        mem_write;
        logic        reg_write;
        logic        csr_we;
    } memory_signals_t;

    // ----- Parameters -----
    localparam REG_WIDTH = $bits(memory_signals_t);

    // ----- Memory pipeline register -----
    memory_signals_t inputs_m;
    memory_signals_t outputs_m;

    assign inputs_m = {
        instr_e_i,
        valid_e_i,
        alu_result_e_i,
        write_data_e_i,
        pc_target_e_i,
        pc_plus4_e_i,
        imm_ext_e_i,
        csr_result_e_i,
        csr_data_e_i,
        csr_addr_e_i,
        rd_e_i,
        width_src_e_i,
        result_src_e_i,
        mem_write_e_i,
        reg_write_e_i,
        csr_we_e_i
    };

    flop #(
        .WIDTH                          (REG_WIDTH)
    ) u_flop_memory_reg (
        // Clock & reset_i
        .clk_i                          (clk_i),
        .reset                          (reset_i),
        .en                             (~stall_m_i),

        // data input
        .D                              (inputs_m),

        // data output
        .Q                              (outputs_m)
    );

    assign {
        instr_m_o,
        valid_m_o,
        alu_result_m_o,
        write_data_m_o,
        pc_target_m_o,
        pc_plus4_m_o,
        imm_ext_m_o,
        csr_result_m_o,
        csr_data_m_o,
        csr_addr_m_o,
        rd_m_o,
        width_src_m_o,
        result_src_m_o,
        mem_write_m_o,
        reg_write_m_o,
        csr_we_m_o
    } = outputs_m;

    // Forwarding mux
    always_comb begin
        case (result_src_m_o)
            `RESULT_ALU:      forward_data_m_o = alu_result_m_o;
            `RESULT_PCTARGET: forward_data_m_o = pc_target_m_o;
            `RESULT_PCPLUS4:  forward_data_m_o = pc_plus4_m_o;
            `RESULT_IMM_EXT:  forward_data_m_o = imm_ext_m_o;
            default:          forward_data_m_o = '0;
        endcase
    end

    reduce u_reduce_width_change (
        // data input
        .BaseResult                     (read_data_m_i),

        // Control input
        .width_src_i                    (width_src_m_o),

        // data output
        .result_o                       (reduced_data_m_o)
    );

endmodule
